module treplo

// Logging levels
pub enum Level {
	panic = 0
	fatal
	error
	warn
	info
	debug
}